** Profile: "SCHEMATIC1-DC op pt"  [ \\gaia.ecs.csus.edu\pheedley\PSpice\examples\eee232\comparator_latching\comparator_latching-PSpiceFiles\SCHEMATIC1\DC op pt.sim ] 

** Creating circuit file "DC op pt.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../comparator_latching-pspicefiles/comparator_latching.lib" 
* From [PSPICE NETLIST] section of t:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.OP
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
