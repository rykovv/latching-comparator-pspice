** Profile: "SCHEMATIC1-testtran"  [ D:\OneDrive\OneDrive - Asian Answers\Documentos\CSUS\EEE232\Projects\Project 1\comparator_latching\comparator_latching-pspicefiles\schematic1\testtran.sim ] 

** Creating circuit file "testtran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../comparator_latching-pspicefiles/comparator_latching.lib" 
* From [PSPICE NETLIST] section of D:\Users\Vladmachine\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN/OP  0 50ns 0 50ps 
.OPTIONS ADVCONV
.OPTIONS ITL4= 100
.OPTIONS RELTOL= 0.0001
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
